class axi_interconnect_wr_ref_model;


endclass
